// -------------------- 7-seg decoder (0..9) --------------------
module sevenseg_decoder (
  parameter bit ACTIVE_LOW = 1   // 1=segments active-low (common anode)
) (
  input  logic [3:0] d,          // BCD 0..9
  output logic [6:0] seg         // a..g
);
  logic [6:0] hi; // active-high
  always_comb unique case (d)
    4'd0: hi=7'b1111110; 4'd1: hi=7'b0110000; 4'd2: hi=7'b1101101; 4'd3: hi=7'b1111001;
    4'd4: hi=7'b0110011; 4'd5: hi=7'b1011011; 4'd6: hi=7'b1011111; 4'd7: hi=7'b1110000;
    4'd8: hi=7'b1111111; 4'd9: hi=7'b1111011; default: hi=7'b0000001; // dash
  endcase
  assign seg = ACTIVE_LOW ? ~hi : hi;
endmodule

// -------------------- Clock ticks --------------------
module pulse_div #(parameter int FCLK=100_000_000, parameter int HZ=1)(
  input  logic clk, rst_n,
  output logic tick
);
  localparam int N = (FCLK/HZ) - 1;
  int c;
  always_ff @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin c<=0; tick<=0; end
    else begin
      tick <= (c==N);
      c    <= (c==N) ? 0 : c+1;
    end
  end
endmodule

// -------------------- Walk timer --------------------
module walk_timer #(
  parameter int WALK_SECS = 10
) (
  input  logic clk, rst_n, tick_1hz, tick_flash,
  input  logic walk_start,             // 1-cycle
  output logic walk_active, walk_done, // pulse on finish
  output logic walk_led,               // flashes while active
  output logic [6:0] secs              // up to 127 secs (we use 0..WALK_SECS)
);
  typedef enum logic {IDLE,RUN} st_t; st_t st;
  logic [6:0] rem; logic led_q;

  always_ff @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin st<=IDLE; rem<=0; walk_done<=0; led_q<=0; end
    else begin
      walk_done <= 0;
      case(st)
        IDLE: if(walk_start) begin st<=RUN; rem<=WALK_SECS; led_q<=0; end
        RUN:  if(tick_1hz) begin
                if(rem==0) begin st<=IDLE; walk_done<=1; end
                else rem <= rem-1;
              end
      endcase
      if(st==RUN && tick_flash) led_q <= ~led_q;
      if(st==IDLE) led_q <= 0;
    end
  end
  assign walk_active = (st==RUN);
  assign walk_led    = led_q;
  assign secs        = rem;
endmodule

// -------------------- Two-digit 7-seg multiplexer --------------------
module sevenseg2 #(
  parameter bit SEG_ACTIVE_LOW = 1,        // segments polarity
  parameter bit AN_ACTIVE_LOW  = 1         // anode/cathode polarity
) (
  input  logic clk, rst_n, tick_mux,
  input  logic [3:0] ones, tens,
  output logic [6:0] seg,
  output logic [3:0] an                    // an[0]=ones, an[1]=tens
);
  logic sel; // 0 ones, 1 tens
  always_ff @(posedge clk or negedge rst_n) begin
    if(!rst_n) sel<=0; else if(tick_mux) sel<=~sel;
  end

  sevenseg_decoder #(.ACTIVE_LOW(SEG_ACTIVE_LOW)) dec(
    .d(sel ? tens : ones), .seg(seg)
  );

  // enable exactly one digit
  always_comb begin
    logic [3:0] hi = sel ? 4'b0010 : 4'b0001;      // active-high intent
    an = AN_ACTIVE_LOW ? ~hi : hi;
  end
endmodule

// -------------------- Top: universal pedestrian display --------------------
module ped_walk_display #(
  parameter int FCLK_HZ       = 100_000_000, // your board clock
  parameter int WALK_SECS     = 10,          // countdown seconds
  parameter int MUX_HZ        = 1000,        // 1–4 kHz typical
  parameter int FLASH_HZ      = 2,           // LED blink rate
  parameter bit SEG_ACTIVE_LOW= 1,           // 1=common-anode segments
  parameter bit AN_ACTIVE_LOW = 1            // 1=common-anode enables
) (
  input  logic clk, rst_n,
  input  logic walk_start,        // pulse from traffic FSM
  output logic walk_done,         // pulse to traffic FSM
  output logic walk_led,          // blink while active
  output logic [6:0] seg,
  output logic [3:0] an
);
  // ticks
  logic t1hz, tmux, tflash;
  pulse_div #(.FCLK(FCLK_HZ), .HZ(1        )) div1 (.clk(clk), .rst_n(rst_n), .tick(t1hz));
  pulse_div #(.FCLK(FCLK_HZ), .HZ(MUX_HZ   )) divm (.clk(clk), .rst_n(rst_n), .tick(tmux));
  pulse_div #(.FCLK(FCLK_HZ), .HZ(2*FLASH_HZ)) divf (.clk(clk), .rst_n(rst_n), .tick(tflash));

  // timer
  logic active; logic [6:0] secs;
  walk_timer #(.WALK_SECS(WALK_SECS)) wt(
    .clk(clk), .rst_n(rst_n), .tick_1hz(t1hz), .tick_flash(tflash),
    .walk_start(walk_start), .walk_active(active), .walk_done(walk_done),
    .walk_led(walk_led), .secs(secs)
  );

  // BCD split
  logic [3:0] ones = secs % 10;
  logic [3:0] tens = (secs/10) % 10;

  // display
  sevenseg2 #(.SEG_ACTIVE_LOW(SEG_ACTIVE_LOW), .AN_ACTIVE_LOW(AN_ACTIVE_LOW)) disp(
    .clk(clk), .rst_n(rst_n), .tick_mux(tmux),
    .ones(ones), .tens(tens), .seg(seg), .an(an)
  );
endmodule
