module clock
(
    input logic counter[5:0],
    input logic PED, 
    input logic mainTraffic[2:0];
    input logic sideTraffic[2:0];
    output logic enable
);

always_comb begin
    enable = 1'b0;
    
        enable = (counter == 6'd15 ||
                  counter == 6'd17 ||
                  counter == 6'd19 ||
                  counter == 6'd27 ||
                  counter == 6'd29);
    end 
end

endmodule
